`define MAX_HOST_NUMBER     32
`define MAX_PLANE_NUMBER    32
`define NO_OF_TAG           1024
