module top
(
    input clk,
    input reset_n,
)

bitmap_manager bitmap_manager(
    .i_clk(clk),
    .i_rst_n(
);
endmodule
